// 





//
