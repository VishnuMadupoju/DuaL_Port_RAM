/* 

   Multi 



*/
